// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
// Created on Sun Oct 26 22:59:03 2025

// synthesis message_off 10175

`timescale 1ns/1ns

module FSM (
    clock,reset,Din,
    Dout);

    input clock;
    input reset;
    input Din;
    tri0 reset;
    tri0 Din;
    output Dout;
    reg Dout;
    reg [5:0] fstate;
    reg [5:0] reg_fstate;
    parameter S0=0,S1=1,S2=2,S3=3,S4=4,S5=5;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or Din)
    begin
        if (reset) begin
            reg_fstate <= S0;
            Dout <= 1'b0;
        end
        else begin
            Dout <= 1'b0;
            case (fstate)
                S0: begin
                    if (~(Din))
                        reg_fstate <= S1;
                    else if (Din)
                        reg_fstate <= S0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S0;

                    Dout <= 1'b0;
                end
                S1: begin
                    if (Din)
                        reg_fstate <= S2;
                    else if (~(Din))
                        reg_fstate <= S1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S1;

                    Dout <= 1'b0;
                end
                S2: begin
                    if (~(Din))
                        reg_fstate <= S3;
                    else if (Din)
                        reg_fstate <= S0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S2;

                    Dout <= 1'b0;
                end
                S3: begin
                    if (Din)
                        reg_fstate <= S4;
                    else if (~(Din))
                        reg_fstate <= S1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S3;

                    Dout <= 1'b0;
                end
                S4: begin
                    if (Din)
                        reg_fstate <= S5;
                    else if (~(Din))
                        reg_fstate <= S3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S4;

                    Dout <= 1'b0;
                end
                S5: begin
                    if (Din)
                        reg_fstate <= S0;
                    else if (~(Din))
                        reg_fstate <= S1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S5;

                    Dout <= 1'b1;
                end
                default: begin
                    Dout <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // FSM
